library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library UART;
use UART.UART_pkg.all;

package UART_tb is
     
end package;
